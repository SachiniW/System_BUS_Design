module char7(c,hEX0);
	input [3:0] c;
	output [6:0] hEX0;
	
	assign hEX0[0] = ((~c[3])&(~c[2])&(~c[1])&(c[0]))|((~c[3])&(c[2])&(~c[1])&(~c[0]))|((c[3])&(~c[2])&(c[1])&(c[0]))|((c[3])&(c[2])&(~c[1])&(c[0]));
	assign hEX0[1] = ((c[2])&(c[1])&(~c[0]))|((c[3])&(c[1])&(c[0]))|((c[3])&(c[2])&(~c[0]))|((~c[3])&(c[2])&(~c[1])&(c[0]));
	assign hEX0[2] = ((~c[3])&(~c[2])&(c[1])&(~c[0]))|((c[3])&(c[2])&(c[1]))|((c[3])&(c[2])&(~c[0]));
	assign hEX0[3] = ((~c[3])&(~c[2])&(~c[1])&(c[0]))|((~c[3])&(c[2])&(~c[1])&(~c[0]))|((c[2])&(c[1])&(c[0]))|((c[3])&(~c[2])&(c[1])&(~c[0]));
	assign hEX0[4] = ((~c[3])&(c[0]))|((~c[3])&(c[2])&(~c[1]))|((c[3])&(~c[2])&(~c[1])&(c[0]));
	assign hEX0[5] = ((c[3])&(c[2])&(~c[1])&(c[0]))|((~c[3])&(~c[2])&(c[0]))|(~(c[3])&(~c[2])&(c[1]))|((~c[3])&(c[1])&(c[0]));
	assign hEX0[6] = ((~c[3])&(~c[2])&(~c[1]))|((~c[3])&(c[2])&(c[1])&(c[0]))|((c[3])&(c[2])&(~c[1])&(~c[0]));
	
endmodule
