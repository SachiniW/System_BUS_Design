module slave_port(
	input clk, 
	input reset,

	input read_en,
	input write_en,

	input master_ready,
	input master_valid,
	
	output reg slave_valid,
	output slave_ready,

	input rx_address,
	input rx_data,

	output slave_tx_done,
	output rx_done,
	output tx_data,


	input [7:0]datain,
	output [11:0]address,
	output [7:0]data,
	
	output read_en_in,
	output reg write_en_in = 0);
	
	
wire slave_ready_IN;
wire slave_ready_OUT;


reg temp2 = 0;
reg temp3 = 0;
reg slave_valid_in = 0;
reg read_en_in1 = 0;
reg write_en_in1 = 0;

assign slave_ready = slave_ready_IN & slave_ready_OUT;
assign read_en_in = rx_done & read_en_in1;
	
slave_in_port SLAVE_IN_PORT(
	.clk(clk), 
	.reset(reset),
	.rx_address(rx_address),
	.rx_data(rx_data),
	.master_valid(master_valid),
	.read_en(read_en),
	.write_en(write_en),
	.slave_ready(slave_ready_IN),
	.rx_done(rx_done),
	.address(address),
	.data(data));
	
slave_out_port SLAVE_OUT_PORT(
	.clk(clk), 
	.reset(reset),
	.master_ready(master_ready),
	.datain(datain),
	.slave_valid(slave_valid),
	.slave_ready(slave_ready_OUT),
	.slave_tx_done(slave_tx_done),
	.tx_data(tx_data));
	

always @ (posedge clk)
begin

	if ((read_en_in1 == 1) & (rx_done == 1) & (slave_valid_in == 0)) 
		slave_valid <= 1;
	else if((slave_tx_done == 1) & (slave_valid_in == 1))
		slave_valid <= 0;
	
	
	if (read_en == 1)
		read_en_in1 <= 1;
	else if (write_en == 1)
	begin
		write_en_in1 <= 1;
		temp2 <= 1;
		temp3 <= 1;
	end

	
	else if ((write_en_in1 == 1) & (rx_done == 1))
		temp2 <= 0;
	else 
	begin
		temp3 <= temp2;
		write_en_in1 <= temp3;
	end
	
	if ((write_en_in1 == 1) & (rx_done == 1))
		write_en_in <= 1;
	if ((write_en_in1 == 0) & (write_en_in == 1))
		write_en_in <= 0;
	if ((rx_done==1) & (read_en_in1 == 1))
		read_en_in1 <= 0;

end
	
endmodule
